Comparador8_inst : Comparador8 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		aeb	 => aeb_sig
	);
