Contador8_inst : Contador8 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
