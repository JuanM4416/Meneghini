Contador16_inst : Contador16 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
