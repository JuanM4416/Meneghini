Registro7_inst : Registro7 PORT MAP (
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		q	 => q_sig,
		shiftout	 => shiftout_sig
	);
