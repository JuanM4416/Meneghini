Comparador7_inst : Comparador7 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		aeb	 => aeb_sig
	);
