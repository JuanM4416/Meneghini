-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Nov 06 15:51:21 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ParteD IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        Q3 : OUT STD_LOGIC;
        Q2 : OUT STD_LOGIC;
        Q1 : OUT STD_LOGIC;
        Q0 : OUT STD_LOGIC
    );
END ParteD;

ARCHITECTURE BEHAVIOR OF ParteD IS
    TYPE type_fstate IS (A,B,E,C,F,D,G);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_Q3 : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x,reg_Q3)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            reg_Q3 <= '0';
            Q3 <= '0';
            Q2 <= '0';
            Q1 <= '0';
            Q0 <= '0';
        ELSE
            reg_Q3 <= '0';
            Q2 <= '0';
            Q1 <= '0';
            Q0 <= '0';
            Q3 <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((x = '0')) THEN
                        reg_fstate <= B;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= G;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    Q0 <= '0';

                    Q1 <= '0';

                    Q2 <= '0';

                    reg_Q3 <= '0';
                WHEN B =>
                    reg_fstate <= C;

                    Q0 <= '0';

                    Q1 <= '1';

                    Q2 <= '1';

                    reg_Q3 <= '0';
                WHEN E =>
                    reg_fstate <= A;

                    Q0 <= '0';

                    Q1 <= '1';

                    Q2 <= '1';

                    reg_Q3 <= '1';
                WHEN C =>
                    IF ((x = '1')) THEN
                        reg_fstate <= E;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= D;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    Q0 <= '1';

                    Q1 <= '1';

                    Q2 <= '1';

                    reg_Q3 <= '1';
                WHEN F =>
                    reg_fstate <= C;

                    Q0 <= '0';

                    Q1 <= '0';

                    Q2 <= '1';

                    reg_Q3 <= '1';
                WHEN D =>
                    reg_fstate <= A;

                    Q0 <= '1';

                    Q1 <= '0';

                    Q2 <= '0';

                    reg_Q3 <= '1';
                WHEN G =>
                    reg_fstate <= F;

                    Q0 <= '0';

                    Q1 <= '0';

                    Q2 <= '0';

                    reg_Q3 <= '1';
                WHEN OTHERS => 
                    reg_Q3 <= 'X';
                    Q2 <= 'X';
                    Q1 <= 'X';
                    Q0 <= 'X';
                    report "Reach undefined state";
            END CASE;
            Q3 <= reg_Q3;
        END IF;
    END PROCESS;
END BEHAVIOR;
